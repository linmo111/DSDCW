//// CORDIC parameters
//`define M  14; // No. of iterations
//`define W  32; // Bit width

// Interface

module CORDIC #(
	parameter M =18,
	parameter W=32

	)(
	input [W-1:0] dataa,
	input clk,
//	input rst,
	input clk_en,
	
	output [W-1:0] result
	);

	// Signals
	reg [W-1:0] x [0:M];
	reg [W-1:0] y [0:M];
	reg [W-1:0] z [0:M]; // Pipeline registers
	reg [M-1:0] di [0:M]; // M-bit direction vector
	reg [W-1:0] e [0:M-1];
//	reg [W-1:0] e [0:M-1] = {
//	 32'b00111111010010010000111111011011,
//	 32'b00111110111011010110001100110001,
//	 32'b00111110011110101101101110110000,
//	 32'b00111101111111001010000110001011,
//	 32'b00111101011111111010101011011110,
//	 
//	 32'b00111100111111111110101010101110,
//	 32'b00111100011111111111101010101010,
//	 32'b00111011111111111111111010101011,
//	 32'b00111011011111111111111110101010,
//	 32'b00111010111111111111111111101111,
//	 
//	 32'b00111010011111111111111111100110,
//	 32'b00111001111111111111111111010101,
//	 32'b00111001011111111111111111010101,
//	 32'b00111000111111111111111111010101,
//	 32'b00111000011111111111111111010101,
//	 
//	 32'b00110111111111111111111011000010,
//	 32'b00110111011111111111110010011100,
//    32'b00110110111111111111110010011100
//
//};
initial begin
	e[0]=32'b00111111010010010000111111011011;
	e[1]=32'b00111110111011010110001100110001;
	e[2]=32'b00111110011110101101101110110000;
	e[3]=32'b00111101111111001010000110001011;
	e[4]=32'b00111101011111111010101011011110;
	
	e[5]=32'b00111100111111111110101010101110;
	e[6]=32'b00111100011111111111101010101010;
	e[7]=32'b00111011111111111111111010101011;
	e[8]=32'b00111011011111111111111110101010;
	e[9]=32'b00111010111111111111111111101111;
	
	e[10]=32'b00111010011111111111111111100110;
	e[11]=32'b00111001111111111111111111010101;
	e[12]=32'b00111001011111111111111111010101;
	e[13]=32'b00111000111111111111111111010101;
	e[14]=32'b00111000011111111111111111010101;
	
	e[15]=32'b00110111111111111111111011000010;
	e[16]=32'b00110111011111111111110010011100;
	e[17]=32'b00110110111111111111110010011100;

	
end

//	assign x[0]=32'b00111111000110110111010011101110;
//	assign y[0]=0;
//	assign z[0] = dataa;
//	assign di = dataa[W-1:W-M]; // MSBs of x



	// CORDIC rotations
	generate
	genvar i;
	for(i=0; i<M; i=i+1) begin : stages
	
		always@ (posedge clk ) begin
		
				if (clk_en) begin
					x[0]=32'b00111111000110110111010011101110;
					y[0]=0;
					z[0] = dataa;
					di[0]=dataa[W-1:W-M];
					x[i+1]=x[i]- ({(di[i]),y[i][30:0]}<<i) ;
					y[i+1]=y[i]+ ({(di[i]),x[i][30:0]}<<i) ;
					z[i+1] =z[i]- ({(di[i]),e[i][30:0]}<<i) ;
					di[i+1]=di[i];
				end
			
		end
		
		
	
	end

	endgenerate

	// Assign output
	assign result = x[M];

	// Initial values

//	assign zi[0] = {1'b1, {(W-1){1'b0}}};

	

endmodule